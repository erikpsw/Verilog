module top_module ( input a, input b, output out );
    
endmodule
