module top_module(
    
    output zero
);// Module body starts after semicolon

endmodule
