module mod_a ( input in1, input in2, output out );
    // Module body
endmodule