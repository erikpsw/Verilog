// synthesis verilog_input_version verilog_2001
module top_module ( 
    input [2:0] sel, 
    input [3:0] data0,
    input [3:0] data1,
    input [3:0] data2,
    input [3:0] data3,
    input [3:0] data4,
    input [3:0] data5,
    output reg [3:0] out   );//

    always@(*) begin  // This is a combinational circuit
        case(sel)
            2'b000:out=data0;
            2'b001:out=data1;
            2'b010:out=data1;
            2'b011:out=data1;
            2'b100:out=data1;
            2'b101:out=data1;
            default:out={4{0}};
        endcase
    end

endmodule
