module top_module ( input a, input b, output out );
    mod_a ins1 (.in1(a),.in1(b),.out(out));
endmodule
