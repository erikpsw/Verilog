module top_module( 
    input a,b,c,
    output w,x,y,z );
    assign w=a,x=b;

endmodule
