module top_module ( input clk, input d, output q );
    my_di
endmodule
