module top_module ( input clk, input d, output q );
    my_dff b1()
endmodule
