module top_module ( input a, input b, output out );
    module top_module ( .out(wc),.in1(wa) );
    endmodule
endmodule
