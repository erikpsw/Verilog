// synthesis verilog_input_version verilog_2001
module top_module (
    input [15:0] scancode,
    output reg left,
    output reg down,
    output reg right,
    output reg up  ); 
    always @(*) begin
        case (scancode)
            16'he06b: 
            default: 
        endcase
    end
endmodule
