module top_module ( input a, input b, output out );
    module top_module ( .out(a),.in1(b),.in2(out) )
endmodule
