module top_module(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);
    a
endmodule
