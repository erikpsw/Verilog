module top_module ( input a, input b, output out );
    mod_a ins1 (.out(a),.in1(b),.in2(out) );
endmodule
