module top_module ( input clk, input d, output q );
    
endmodule
