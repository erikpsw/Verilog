module top_module ( input a, input b, output out );
    mod_a instance1 ( wa, wb, wc );
endmodule