module top_module ( input a, input b, output out );
    module top_module ( input a, input b, output out );
    endmodule
endmodule
